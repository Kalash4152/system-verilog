// AND gate module
module and_gate(
    input a,
    input b,
    output y
);
    assign y = a & b;  // AND operation
endmodule
